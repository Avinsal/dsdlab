module Q1(a,b,c,d,En,f);
input a,b,c,d;
input En;
output f;
output z;
wire [0:15]y;
wire [0:3]w;
assign w={a,b,c,d};
dec4to16 s1(w,y,En);
assign f=y[1]|y[3]|y[6]|y[7]|y[9]|y[14]|y[15];
endmodule

module dec4to16(w,y,En);
input [0:3]w;
input En;
output [0:15]y;
reg [0:15]y;
always@(w or En)
begin 
if(En==0)
y=16'b0000000000000000;
else
case(w)
0:y=16'b1000000000000000;
1:y=16'b0100000000000000;
2:y=16'b0010000000000000;
3:y=16'b0001000000000000;
4:y=16'b0000100000000000;
5:y=16'b0000010000000000;
6:y=16'b0000001000000000;
7:y=16'b0000000100000000;
8:y=16'b0000000010000000;
9:y=16'b0000000001000000;
10:y=16'b0000000000100000;
11:y=16'b0000000000010000;
12:y=16'b0000000000001000;
13:y=16'b0000000000000100;
14:y=16'b0000000000000010;
15:y=16'b0000000000000001;
endcase
end
endmodule





